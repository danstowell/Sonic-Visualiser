BZh91AY&SYē�� m_�ryc���o߰����`�=�s���{ �@����@ ���3T�"h�M4h  � �h� h �U�L   ���5D���� �#`�M4"jjOBM�h�G��P���z�� �@ᦙ�&�`L#��i���
�@@C��0MF�bbi���i�0HC�|��� �~J%��$M"!uI-�}�"I||�����GVG�����G��Ơ�2 ~����m���Ya�'��T��A��u�,����̪?��]��U�)=ޯ_{OWυ��͓��6hW�F7�A �O'N���U{t9-��z�쭃��F���PD�i�>o���Z�Ƹ�|�|���AEB����A�P��A�J6���>���Ӎ8�*�<�2m��%В���DN\2�*��@5��mjn���d!��2������˶S%�D���j`�MCFO��:y�����s35��_S�z3�s`�6�.2F�(�K�q��Qr.E�9hΩŐ           � ���kj%�t��ȉEm����R�� �%  +7+��P�$���m�+��2) X�	m����`�c��  
�TYH����.�ck?����a#5���B:c��6$>����zL�s�9�@�>S�Ø`�������8L���8�)�ʗR���v��V�RH$K�-(�D#� �H) � \u�lm�a梮�M��WS.6��m�}k�@�U $	T���z��Lj7�h�ʜ�I_I^0�Ê}oZ� $�&s�&���Q2�*n�t�ƚX֔��G.�c�/l�"��[1Qq����3{u!i���ժ)PlW��
@m2[�*���M���v�u�
��;3*���f2;��p^.�N!�5�G@�n�0�y1�-�
��jB����
�R=���x�
�E��P�N�0��%� �F���Z���R�E�TYU xeyU���p�Ņ�a(���hQ�������({����R���(��w�i�O�Y�U��U�8���Q���O�3��)!�e|�W����<	���R��6	�A�f̺m��� :А���(��b�3��{��9��B��oɳ�G�P���+u�1ӬV�{ie­%XJ*�JH(���pہ���r8������)
i�]�𤊺���?��|��qq����f�(�e*��3��5 �Z��;H�5�a�EJ����^�r8�����({��'v�vX���y�y�O������uh��"���E����ɸ��{����h����3�V��6XhM�ӛ��m�8��)�0ٲ*���k�����I%�Ѵ{*'�����x HB(��
6�85�a�Mo\&�t�t(
��A\����KT����7��,{@�<`�<E{wm�mNŘ�_g�>�ӹ6i�v";Ӑ�狃oE��μZ��S�k���U���k��n�9���s�%Y��Z��f��y�~x�W�|�1�7�J�i���/��P4ܽC,Ųձehw��b�ge6�8�0*���3�/=l4�AcohT88�\�NN�vg*�]mwheXWH�ͮZ���79�!���:I�e����865yY����}
'FUL����-���+��pv���Cܛ�Ut�f���/p*�-�¢� H"!&��M=��4*��P���5;$�Z�Sl�A��+2\.l�tx��\��L8:,m�̴�_4�gƷh��)
���9L���l��/Ք/V��gW����A؎ˡl�f.c�n�h�#�1�4YU�
7N����E�#'qk��sUfzyoGn����ܴu�I�'m�eg	�-�����á��}g�;�p ��P
�(�`۬�ՉWr=Z`�Y��̬O�zG..��7r�/_�x5�L*О��7*�ݒ�����~h��f\����fR6�b*�k,����*Ttu\\b�����*W�ž�']�7��A�h�0"8��UVc���@�W�ыC��5������j�C�;c�k�6>�n���p�|���d�\r-%R�j<j��VgL�Wt8����Ѥ	*I$�H���@,�=&� �%�ɓ��0��&x�1�h$��/��sYR9*��in(�*ܐ��/EC�	&`%��d�T ��5��L)e!J0��(DśX��&	����H����C��%�Y�	.wȨ�q��T�N~ʽ�E����k�Yq���� K�c;�;g��T	 Bo)�u�y��<��	a�a���|̡v���轖��բ�3�x���r��8�K:oz�7y�:�����K:"��ꪙ���,���#�$��e>2��"��^;��6�nt����SW�N�I�-/�cs���#�`+��6�����1x7)�(��_"���E�ն��O�T�b�qmuKF���6w`��)�&���b1;���=B�?�������b/���0i��t����nz��(`��ɚ?#�}���=��0��W����٫ּ�0ka6*�ؽ��l�yi� �*q� ��8H�n��T��ߌ�-��6b1�*22I�X�dFEdD�da�@i���/!��t1��Hw��'�	��08�r���@ȴ��-�c��Ϸ|�87�V+${��^���l�	�v��ёח���o0l3Of�j=�>��>�z=�<>Ȣ�j���d]=�^Z��#�,ږ˜}��h�]m�ڲf�����l��`��ww7a���SK��1[l���q��u��'�7�i��Ю�	���II\Z��IT�����y�_��(�T����0�I �| s>����'�%duk�|.W���X�5��ϱ�(���f^��#̩$��Q���mXܩA��	mi�4)��1P ��)�߸ڻ"}A@]Q�RU��ha!�F��L�'dT[;/_&%�R]c�L�IE��A^.�����B�:�HuBYv���RK����y]������j��~�/�ͱt�S�76޴S���G7G3�x)N�b��q�])S����C5�����@����7C|�MqIH�:��O Zyo�%/\y���|m4ҹ`���v�����̤i��vY**)��+��Ş�^��M��1vI��+5���c��!�F������|d+.)�d����_^�@ͳ�st���K��8�EɆ6L/.��k�י��p#'Z�J]ݥy���&�%���t/4���/ތ6��"�%I4w�ǐ_�4�ZIҧ����h�46�j���:N�c���LL���3�1Ύ���c��nU�N��O��:�~�����H�
�|~@